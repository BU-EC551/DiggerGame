`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:47:45 03/23/2015 
// Design Name: 
// Module Name:    vgacontroller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vgacontroller(clk100m, clk40m,
							hs, vs, 
							r0, r1, r2, r3, 
							g0, g1, g2, g3,
							b0, b1, b2, b3,
							dig_posx,
							dig_posy,
							gob_posx,
							gob_posy,
							dmov, gmov,
					      vgaram_we,
					      vgaram_addra,
					      vgaram_dina,
					      vgaram_douta,	
							score,
							game_over,
							mb0_exist,
							mb1_exist,
							mb2_exist,
							mb3_exist,
							mb4_exist
							);
							
   input      clk100m;
	input      clk40m;
	input  [2:0] dmov;
	input  [2:0] gmov;
	
	input    	 vgaram_we;
	input [7:0]	 vgaram_addra;
	input [3:0]	 vgaram_dina;
	input wire [9:0]  score;
	input        game_over;
	input [1:0] mb0_exist;
	input [1:0] mb1_exist;
	input [1:0] mb2_exist;
	input [1:0] mb3_exist;
	input [1:0] mb4_exist;
	output [3:0]  vgaram_douta;
	
   output     hs;
   output     vs;
	//12-bit rgb
   output     r0;
   output     r1;
   output     r2;
   output     r3;
   output     g0;
   output     g1;
   output     g2;
   output     g3;
   output     b0;
   output     b1;
   output     b2;
   output     b3;
   
	output	[9:0]	dig_posx;
	output	[9:0]	dig_posy;
	output	[9:0]	gob_posx;
	output 	[9:0]	gob_posy;
	
   wire       clk25m;
   wire       clk1hz;
   wire       clk100hz;
	wire       clk5m;

   wire [10:0] vcnt;
   wire [10:0] hcnt;
   wire       ven;
   wire       hen;
	
   wire [11:0] colors;
   wire [5:0] colors3;

   assign {r3, r2, r1, r0, g3, g2, g1, g0, b3, b2, b1, b0} = colors;
	
	 
	 
	clock clock_port_map(.clk50m(clk100m), 
	                     .clk25m(clk25m), 
								.clk100hz(clk100hz), 
								.clk1hz(clk1hz), 
								.clk5m(clk5m)
								);
   
   
   pixelcnt pixelcnt_port_map(.clk25m(clk40m), 
	                           .hcntout(hcnt), 
										.vcntout(vcnt)
										);
   
   
   vgasig vgasig_port_map(.clk25m(clk40m), 
	                       .hcnt(hcnt), 
								  .vcnt(vcnt), 
								  .hsync(hs), 
								  .vsync(vs), 
								  .henable(hen), 
								  .venable(ven)
								  );
   
   
   vgacolor vgacolor_port_map(.clk5m(clk5m), .clk100m(clk100m), .clk25m(clk40m), .clk100hz(clk100hz),
										.clk_vgaram(clk100m), .vgaram_we(vgaram_we), 
										.vgaram_addra(vgaram_addra), 
										.vgaram_dina(vgaram_dina), .vgaram_douta(vgaram_douta),
										
	                           .hen(hen), .ven(ven), .hpos(hcnt), .vpos(vcnt),
										.dmov(dmov), .gmov(gmov), 
										.colors(colors),
										.dig_posx(dig_posx),
										.dig_posy(dig_posy),
										.gob_posx(gob_posx),
										.gob_posy(gob_posy),
										.score(score),
										.game_over(game_over),
										.mb0_exist(mb0_exist),
										 .mb1_exist(mb1_exist),
										 .mb2_exist(mb2_exist),
										 .mb3_exist(mb3_exist),
										 .mb4_exist(mb4_exist)
										);
   
endmodule


