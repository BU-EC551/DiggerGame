`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:58:49 03/21/2015 
// Design Name: 
// Module Name:    map 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module map(Clk,rst,Digx,Digy,Gobx,Goby, out,up,down,left,right,value
    );
	input Clk,rst;
	input [3:0] Digx,Digy,Gobx,Goby;
	input [2:0] value;	//save for money bag
	output [2:0] out;
	output [2:0] up,down,left,right;
	wire [3:0] xup,yup,xdown,ydown,xleft,yleft,xright,yright;
	 reg [3:0] xbdy,ybdy;
	 initial xbdy=4'd10;
	 initial ybdy=4'd15;
	reg [2:0] memory [0:10][0:15];
	
	initial begin
		memory[0][0]=3'd0;
		memory[0][1]=3'd3;
		memory[0][2]=3'd3;
		memory[0][3]=3'd3;
		memory[0][4]=3'd5;
		memory[0][5]=3'd3;
		memory[0][6]=3'd3;
		memory[0][7]=3'd3;
		memory[0][8]=3'd3;
		memory[0][9]=3'd3;
		memory[0][10]=3'd0;
		memory[0][11]=3'd0;
		memory[0][12]=3'd0;
		memory[0][13]=3'd0;
		memory[0][14]=3'd0;
		memory[1][0]=3'd0;
		memory[1][1]=3'd3;
		memory[1][2]=3'd3;
		memory[1][3]=3'd4;
		memory[1][4]=3'd4;
		memory[1][5]=3'd3;
		memory[1][6]=3'd3;
		memory[1][7]=3'd4;
		memory[1][8]=3'd3;
		memory[1][9]=3'd3;
		memory[1][10]=3'd0;
		memory[1][11]=3'd3;
		memory[1][12]=3'd5;
		memory[1][13]=3'd3;
		memory[1][14]=3'd3;
		memory[2][0]=3'd0;
		memory[2][1]=3'd5;
		memory[2][2]=3'd3;
		memory[2][3]=3'd4;
		memory[2][4]=3'd4;
		memory[2][5]=3'd3;
		memory[2][6]=3'd3;
		memory[2][7]=3'd4;
		memory[2][8]=3'd3;
		memory[2][9]=3'd3;
		memory[2][10]=3'd0;
		memory[2][11]=3'd3;
		memory[2][12]=3'd3;
		memory[2][13]=3'd3;
		memory[2][14]=3'd3;
		memory[3][0]=3'd0;
		memory[3][1]=3'd3;
		memory[3][2]=3'd3;
		memory[3][3]=3'd4;
		memory[3][4]=3'd4;
		memory[3][5]=3'd5;
		memory[3][6]=3'd3;
		memory[3][7]=3'd3;
		memory[3][8]=3'd3;
		memory[3][9]=3'd3;
		memory[3][10]=3'd0;
		memory[3][11]=3'd3;
		memory[3][12]=3'd4;
		memory[3][13]=3'd4;
		memory[3][14]=3'd4;
		memory[4][0]=3'd0;
		memory[4][1]=3'd3;
		memory[4][2]=3'd3;
		memory[4][3]=3'd4;
		memory[4][4]=3'd4;
		memory[4][5]=3'd3;
		memory[4][6]=3'd3;
		memory[4][7]=3'd4;
		memory[4][8]=3'd3;
		memory[4][9]=3'd3;
		memory[4][10]=3'd0;
		memory[4][11]=3'd3;
		memory[4][12]=3'd4;
		memory[4][13]=3'd4;
		memory[4][14]=3'd4;
		memory[5][0]=3'd0;
		memory[5][1]=3'd0;
		memory[5][2]=3'd3;
		memory[5][3]=3'd4;
		memory[5][4]=3'd4;
		memory[5][5]=3'd3;
		memory[5][6]=3'd3;
		memory[5][7]=3'd4;
		memory[5][8]=3'd3;
		memory[5][9]=3'd3;
		memory[5][10]=3'd0;
		memory[5][11]=3'd3;
		memory[5][12]=3'd3;
		memory[5][13]=3'd3;
		memory[5][14]=3'd3;
		memory[6][0]=3'd3;
		memory[6][1]=3'd0;
		memory[6][2]=3'd3;
		memory[6][3]=3'd3;
		memory[6][4]=3'd3;
		memory[6][5]=3'd3;
		memory[6][6]=3'd5;
		memory[6][7]=3'd0;
		memory[6][8]=3'd5;
		memory[6][9]=3'd3;
		memory[6][10]=3'd0;
		memory[6][11]=3'd3;
		memory[6][12]=3'd3;
		memory[6][13]=3'd3;
		memory[6][14]=3'd3;
		memory[7][0]=3'd3;
		memory[7][1]=3'd0;
		memory[7][2]=3'd0;
		memory[7][3]=3'd0;
		memory[7][4]=3'd0;
		memory[7][5]=3'd3;
		memory[7][6]=3'd3;
		memory[7][7]=3'd0;
		memory[7][8]=3'd3;
		memory[7][9]=3'd3;
		memory[7][10]=3'd0;
		memory[7][11]=3'd3;
		memory[7][12]=3'd3;
		memory[7][13]=3'd3;
		memory[7][14]=3'd3;
		memory[8][0]=3'd4;
		memory[8][1]=3'd3;
		memory[8][2]=3'd3;
		memory[8][3]=3'd3;
		memory[8][4]=3'd0;
		memory[8][5]=3'd3;
		memory[8][6]=3'd3;
		memory[8][7]=3'd0;
		memory[8][8]=3'd3;
		memory[8][9]=3'd3;
		memory[8][10]=3'd0;
		memory[8][11]=3'd3;
		memory[8][12]=3'd3;
		memory[8][13]=3'd3;
		memory[8][14]=3'd4;
		memory[9][0]=3'd4;
		memory[9][1]=3'd4;
		memory[9][2]=3'd3;
		memory[9][3]=3'd3;
		memory[9][4]=3'd0;
		memory[9][5]=3'd0;
		memory[9][6]=3'd0;
		memory[9][7]=3'd0;
		memory[9][8]=3'd0;
		memory[9][9]=3'd0;
		memory[9][10]=3'd0;
		memory[9][11]=3'd3;
		memory[9][12]=3'd3;
		memory[9][13]=3'd4;
		memory[9][14]=3'd4;
	//boundary	
		memory[10][0]=3'd7;
		memory[10][1]=3'd7;
		memory[10][2]=3'd7;
		memory[10][3]=3'd7;
		memory[10][4]=3'd7;
		memory[10][5]=3'd7;
		memory[10][6]=3'd7;
		memory[10][7]=3'd7;
		memory[10][8]=3'd7;
		memory[10][9]=3'd7;
		memory[10][10]=3'd7;
		memory[10][11]=3'd7;
		memory[10][12]=3'd7;
		memory[10][13]=3'd7;
		memory[10][14]=3'd7;	
		memory[0][15]=3'd7;
		memory[1][15]=3'd7;
		memory[2][15]=3'd7;
		memory[3][15]=3'd7;
		memory[4][15]=3'd7;
		memory[5][15]=3'd7;
		memory[6][15]=3'd7;
		memory[7][15]=3'd7;
		memory[8][15]=3'd7;
		memory[9][15]=3'd7;
		memory[10][15]=3'd7;
	end
	
	assign out=memory[Digx][Digy];
	assign 	xup=(Gobx>0)? Gobx-1 :xbdy;
	assign	yup=Goby;
	assign	xdown=(Gobx<9)?Gobx+1:xbdy;
	assign	ydown=Goby;
	assign	xleft=Gobx;
	assign	yleft=(Goby>0)?Goby-1:ybdy;
	assign	xright=Gobx;
	assign	yright=(Goby<14)?Goby+1:ybdy;	
	assign up=memory[xup][yup];
	assign down=memory[xdown][ydown];
	assign left=memory[xleft][yleft];
	assign right=memory[right][yright];
	
	always @(negedge Clk) begin
		if (rst) begin
		memory[0][0]<=3'd0;
		memory[0][1]<=3'd3;
		memory[0][2]<=3'd3;
		memory[0][3]<=3'd3;
		memory[0][4]<=3'd5;
		memory[0][5]<=3'd3;
		memory[0][6]<=3'd3;
		memory[0][7]<=3'd3;
		memory[0][8]<=3'd3;
		memory[0][9]<=3'd3;
		memory[0][10]<=3'd0;
		memory[0][11]<=3'd0;
		memory[0][12]<=3'd0;
		memory[0][13]<=3'd0;
		memory[0][14]<=3'd0;
		memory[1][0]<=3'd0;
		memory[1][1]<=3'd3;
		memory[1][2]<=3'd3;
		memory[1][3]<=3'd4;
		memory[1][4]<=3'd4;
		memory[1][5]<=3'd3;
		memory[1][6]<=3'd3;
		memory[1][7]<=3'd4;
		memory[1][8]<=3'd3;
		memory[1][9]<=3'd3;
		memory[1][10]<=3'd0;
		memory[1][11]<=3'd3;
		memory[1][12]<=3'd5;
		memory[1][13]<=3'd3;
		memory[1][14]<=3'd3;
		memory[2][0]<=3'd0;
		memory[2][1]<=3'd5;
		memory[2][2]<=3'd3;
		memory[2][3]<=3'd4;
		memory[2][4]<=3'd4;
		memory[2][5]<=3'd3;
		memory[2][6]<=3'd3;
		memory[2][7]<=3'd4;
		memory[2][8]<=3'd3;
		memory[2][9]<=3'd3;
		memory[2][10]<=3'd0;
		memory[2][11]<=3'd3;
		memory[2][12]<=3'd3;
		memory[2][13]<=3'd3;
		memory[2][14]<=3'd3;
		memory[3][0]<=3'd0;
		memory[3][1]<=3'd3;
		memory[3][2]<=3'd3;
		memory[3][3]<=3'd4;
		memory[3][4]<=3'd4;
		memory[3][5]<=3'd5;
		memory[3][6]<=3'd3;
		memory[3][7]<=3'd3;
		memory[3][8]<=3'd3;
		memory[3][9]<=3'd3;
		memory[3][10]<=3'd0;
		memory[3][11]<=3'd3;
		memory[3][12]<=3'd4;
		memory[3][13]<=3'd4;
		memory[3][14]<=3'd4;
		memory[4][0]<=3'd0;
		memory[4][1]<=3'd3;
		memory[4][2]<=3'd3;
		memory[4][3]<=3'd4;
		memory[4][4]<=3'd4;
		memory[4][5]<=3'd3;
		memory[4][6]<=3'd3;
		memory[4][7]<=3'd4;
		memory[4][8]<=3'd3;
		memory[4][9]<=3'd3;
		memory[4][10]<=3'd0;
		memory[4][11]<=3'd3;
		memory[4][12]<=3'd4;
		memory[4][13]<=3'd4;
		memory[4][14]<=3'd4;
		memory[5][0]<=3'd0;
		memory[5][1]<=3'd0;
		memory[5][2]<=3'd3;
		memory[5][3]<=3'd4;
		memory[5][4]<=3'd4;
		memory[5][5]<=3'd3;
		memory[5][6]<=3'd3;
		memory[5][7]<=3'd4;
		memory[5][8]<=3'd3;
		memory[5][9]<=3'd3;
		memory[5][10]<=3'd0;
		memory[5][11]<=3'd3;
		memory[5][12]<=3'd3;
		memory[5][13]<=3'd3;
		memory[5][14]<=3'd3;
		memory[6][0]<=3'd3;
		memory[6][1]<=3'd0;
		memory[6][2]<=3'd3;
		memory[6][3]<=3'd3;
		memory[6][4]<=3'd3;
		memory[6][5]<=3'd3;
		memory[6][6]<=3'd5;
		memory[6][7]<=3'd0;
		memory[6][8]<=3'd5;
		memory[6][9]<=3'd3;
		memory[6][10]<=3'd0;
		memory[6][11]<=3'd3;
		memory[6][12]<=3'd3;
		memory[6][13]<=3'd3;
		memory[6][14]<=3'd3;
		memory[7][0]<=3'd3;
		memory[7][1]<=3'd0;
		memory[7][2]<=3'd0;
		memory[7][3]<=3'd0;
		memory[7][4]<=3'd0;
		memory[7][5]<=3'd3;
		memory[7][6]<=3'd3;
		memory[7][7]<=3'd0;
		memory[7][8]<=3'd3;
		memory[7][9]<=3'd3;
		memory[7][10]<=3'd0;
		memory[7][11]<=3'd3;
		memory[7][12]<=3'd3;
		memory[7][13]<=3'd3;
		memory[7][14]<=3'd3;
		memory[8][0]<=3'd4;
		memory[8][1]<=3'd3;
		memory[8][2]<=3'd3;
		memory[8][3]<=3'd3;
		memory[8][4]<=3'd0;
		memory[8][5]<=3'd3;
		memory[8][6]<=3'd3;
		memory[8][7]<=3'd0;
		memory[8][8]<=3'd3;
		memory[8][9]<=3'd3;
		memory[8][10]<=3'd0;
		memory[8][11]<=3'd3;
		memory[8][12]<=3'd3;
		memory[8][13]<=3'd3;
		memory[8][14]<=3'd4;
		memory[9][0]<=3'd4;
		memory[9][1]<=3'd4;
		memory[9][2]<=3'd3;
		memory[9][3]<=3'd3;
		memory[9][4]<=3'd0;
		memory[9][5]<=3'd0;
		memory[9][6]<=3'd0;
		memory[9][7]<=3'd0;
		memory[9][8]<=3'd0;
		memory[9][9]<=3'd0;
		memory[9][10]<=3'd0;
		memory[9][11]<=3'd3;
		memory[9][12]<=3'd3;
		memory[9][13]<=3'd4;
		memory[9][14]<=3'd4;

		end else memory[Digx][Digy]<=3'd0;
	end

endmodule

