`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:06:40 03/25/2015 
// Design Name: 
// Module Name:    keyboardtest 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module keyboardtest( 
	input wire clk, // Clock pin form keyboard 
	input wire data, //Data pin form keyboard 
	output reg [7:0] key_out, //Printing input data to key_out
	output reg sample //the posedge of sample denote the key_out is a valid screen output
	); 
	reg [7:0] data_curr; 
	reg [7:0] data_pre; 
	reg [3:0] b; 
	reg flag; 
 
	initial 
		begin 
		b<=4'h1; 
		flag<=1'b0; 
		data_curr<=8'hf0; 
		data_pre<=8'hf0; 
		key_out<=8'hf0;
		end 
 
	always @(negedge clk) //Activating at negative edge of clock from keyboard 
	
	begin 
 
	case(b) 
	1:; //first bit 
	2:data_curr[0]<=data; 
	3:data_curr[1]<=data; 
	4:data_curr[2]<=data; 
	5:data_curr[3]<=data; 
	6:data_curr[4]<=data; 
	7:data_curr[5]<=data; 
	8:data_curr[6]<=data; 
	9:data_curr[7]<=data; 
	10:flag<=1'b1; //Parity bit 
	11:flag<=1'b0; //Ending bit 
 
	endcase 
 
	if(b<=10) 
	b<=b+1; 
 
	else if(b==11) 
	b<=1; 
 
 
	end 
 
	always@(posedge flag) // Printing data obtained to led 
	begin 
 
	 if(data_curr==8'hf0 && data_pre!=8'h58)begin //capslock do not generate any output
	   key_out<=data_pre;
	   sample <= 1; end
	 else begin
	   data_pre<=data_curr;
	   sample <=0; end
	end 
	
	

endmodule


